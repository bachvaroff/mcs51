// XAPP052

module LFSR (CLK, E, RESET, SEED_VAL, LFSR_VAL);

parameter NUM_BITS = 32;

input wire CLK;
input wire E;
input wire RESET;
input wire [(NUM_BITS - 1):0] SEED_VAL;
output wire [(NUM_BITS - 1):0] LFSR_VAL;

reg [NUM_BITS:1] LFSR;
wire XNOR;

assign LFSR_VAL = LFSR;

generate
	case (NUM_BITS)
		3: assign XNOR = LFSR[3] ^ ~LFSR[2];
		4: assign XNOR = LFSR[4] ^ ~LFSR[3];
		5: assign XNOR = LFSR[5] ^ ~LFSR[3];
		6: assign XNOR = LFSR[6] ^ ~LFSR[5];
		7: assign XNOR = LFSR[7] ^ ~LFSR[6];
		8: assign XNOR = LFSR[8] ^ ~LFSR[6] ^ ~LFSR[5] ^ ~LFSR[4];
		9: assign XNOR = LFSR[9] ^ ~LFSR[5];
		10: assign XNOR = LFSR[10] ^ ~LFSR[7];
		11: assign XNOR = LFSR[11] ^ ~LFSR[9];
		12: assign XNOR = LFSR[12] ^ ~LFSR[6] ^ ~LFSR[4] ^ ~LFSR[1];
		13: assign XNOR = LFSR[13] ^ ~LFSR[4] ^ ~LFSR[3] ^ ~LFSR[1];
		14: assign XNOR = LFSR[14] ^ ~LFSR[5] ^ ~LFSR[3] ^ ~LFSR[1];
		15: assign XNOR = LFSR[15] ^ ~LFSR[14];
		16: assign XNOR = LFSR[16] ^ ~LFSR[15] ^ ~LFSR[13] ^ ~LFSR[4];
		17: assign XNOR = LFSR[17] ^ ~LFSR[14];
		18: assign XNOR = LFSR[18] ^ ~LFSR[11];
		19: assign XNOR = LFSR[19] ^ ~LFSR[6] ^ ~LFSR[2] ^ ~LFSR[1];
		20: assign XNOR = LFSR[20] ^ ~LFSR[17];
		21: assign XNOR = LFSR[21] ^ ~LFSR[19];
		22: assign XNOR = LFSR[22] ^ ~LFSR[21];
		23: assign XNOR = LFSR[23] ^ ~LFSR[18];
		24: assign XNOR = LFSR[24] ^ ~LFSR[23] ^ ~LFSR[22] ^ ~LFSR[17];
		25: assign XNOR = LFSR[25] ^ ~LFSR[22];
		26: assign XNOR = LFSR[26] ^ ~LFSR[6] ^ ~LFSR[2] ^ ~LFSR[1];
		27: assign XNOR = LFSR[27] ^ ~LFSR[5] ^ ~LFSR[2] ^ ~LFSR[1];
		28: assign XNOR = LFSR[28] ^ ~LFSR[25];
		29: assign XNOR = LFSR[29] ^ ~LFSR[27];
		30: assign XNOR = LFSR[30] ^ ~LFSR[6] ^ ~LFSR[4] ^ ~LFSR[1];
		31: assign XNOR = LFSR[31] ^ ~LFSR[28];
		32: assign XNOR = LFSR[32] ^ ~LFSR[22] ^ ~LFSR[2] ^ ~LFSR[1];
		64: assign XNOR = LFSR[64] ^ ~LFSR[63] ^ ~LFSR[61] ^ ~LFSR[60];
	endcase
endgenerate

always @(posedge CLK) begin
	if (E) begin
		if (RESET) LFSR <= SEED_VAL;
		else LFSR <= { LFSR[(NUM_BITS - 1):1], XNOR };
	end;
end

endmodule
