module decode_8seg(OE, tetrade, dot, leds_val);

input wire OE;
input wire [3:0] tetrade;
input wire dot;
output wire [7:0] leds_val; /* { dot, g, f, e, d, c, b, a } */

reg [7:0] leds;

assign leds_val = leds;

always @(*) begin
	if (!OE) begin
		leds <= 8'b00000000;
	end else begin
		case (tetrade)
			4'b0000: leds <= { dot, 7'b0111111 }; /* 0. */
			4'b0001: leds <= { dot, 7'b0000110 }; /* 1. */
			4'b0010: leds <= { dot, 7'b1011011 }; /* 2. */
			4'b0011: leds <= { dot, 7'b1001111 }; /* 3. */
			4'b0100: leds <= { dot, 7'b1100110 }; /* 4. */
			4'b0101: leds <= { dot, 7'b1101101 }; /* 5. */
			4'b0110: leds <= { dot, 7'b1111101 }; /* 6. */
			4'b0111: leds <= { dot, 7'b0000111 }; /* 7. */
			4'b1000: leds <= { dot, 7'b1111111 }; /* 8. */
			4'b1001: leds <= { dot, 7'b1101111 }; /* 9. */
			4'b1010: leds <= { dot, 7'b1110111 }; /* A. */
			4'b1011: leds <= { dot, 7'b1111100 }; /* b. */
			4'b1100: leds <= { dot, 7'b0111001 }; /* C. */
			4'b1101: leds <= { dot, 7'b1011110 }; /* d. */
			4'b1110: leds <= { dot, 7'b1111001 }; /* E. */
			4'b1111: leds <= { dot, 7'b1110001 }; /* F. */
		endcase
	end
end

endmodule

